module spi_regs (
	input sck,
	input mosi,
	output reg miso,
	input csn,
	
	output [127:0] data
);

	
endmodule